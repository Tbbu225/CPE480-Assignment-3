


module tacky_processor(halt, reset, clk);

endmodule
